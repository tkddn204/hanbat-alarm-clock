






// DIGITAL_CLOCK.v

module DIGITAL_CLOCK(
	RESETN, CLK,
	KEY,
   LCD_E, LCD_RS, LCD_RW,
	LCD_DATA, PIEZO
);

input RESETN, CLK;
input [4:0] KEY;
output wire LCD_E, LCD_RS, LCD_RW, PIEZO;
output wire [7:0] LCD_DATA;

wire MERIDIAN;
wire [16:0] ALARM_TIME;
wire [16:0] CURRENT_TIME;
wire [15:0] CURRENT_DATE;

wire [16:0] SETTING_ALARM_TIME;
wire [16:0] SETTING_CURRENT_TIME;
wire [15:0] SETTING_CURRENT_DATE;

wire [7:0] CURRENT_H10, CURRENT_H1, CURRENT_M10, CURRENT_M1, CURRENT_S10, CURRENT_S1;
wire [7:0] CURRENT_Y10, CURRENT_Y1, CURRENT_MT10, CURRENT_MT1, CURRENT_D10, CURRENT_D1;
wire [7:0] ALARM_H10, ALARM_H1, ALARM_M10, ALARM_M1, ALARM_S10, ALARM_S1;

wire [5:0] MODE;
wire SETTING, ALARM_SETTING, SETTING_OK;

wire ALARM_ENABLE, ALARM_DOING;

// Key Controller
KEY_CONT key_cont(
	RESETN, CLK,
	KEY, CURRENT_TIME, CURRENT_DATE, ALARM_TIME,
	MODE, ALARM_ENABLE, SETTING, ALARM_SETTING, SETTING_OK,
	SETTING_CURRENT_TIME, SETTING_CURRENT_DATE, SETTING_ALARM_TIME, MERIDIAN
);

// Time Calculator
TIME_CAL time_cal(
	RESETN, CLK,
	SETTING_CURRENT_TIME, SETTING_CURRENT_DATE, SETTING_ALARM_TIME,
	MODE[0], MODE[5], SETTING, ALARM_SETTING, SETTING_OK,
	CURRENT_TIME, CURRENT_DATE, ALARM_TIME,
);

// (current time) and (alarm time) compare
TIME_COMPARE time_compare(
	RESETN, CLK,
	ALARM_ENABLE, CURRENT_TIME, ALARM_TIME,
	ALARM_DOING
);

// PIEZO
PIEZO_UNIT piezo_unit(
	RESETN, CLK,
	ALARM_ENABLE, ALARM_DOING,
	PIEZO
);

// DISPLAY decoder
DISPLAY_DECODER display_decoder(
	RESETN, CLK,
	CURRENT_TIME, CURRENT_DATE, ALARM_TIME,
	CURRENT_H10, CURRENT_H1, CURRENT_M10, CURRENT_M1, CURRENT_S10, CURRENT_S1,
	CURRENT_Y10, CURRENT_Y1, CURRENT_MT10, CURRENT_MT1, CURRENT_D10, CURRENT_D1,
	ALARM_H10, ALARM_H1, ALARM_M10, ALARM_M1, ALARM_S10, ALARM_S1
);

/// DISPLAY Controller
DISPLAY_CONT display_cont(
	RESETN, CLK,
	CURRENT_H10, CURRENT_H1, CURRENT_M10, CURRENT_M1, CURRENT_S10, CURRENT_S1, MERIDIAN,
	CURRENT_Y10, CURRENT_Y1, CURRENT_MT10, CURRENT_MT1, CURRENT_D10, CURRENT_D1,
	ALARM_H10, ALARM_H1, ALARM_M10, ALARM_M1, ALARM_S10, ALARM_S1,
	MODE, ALARM_ENABLE, ALARM_DOING,
	LCD_E, LCD_RS, LCD_RW,
	LCD_DATA
);

endmodule
