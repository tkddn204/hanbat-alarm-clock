






// DIGITAL_CLOCK.v

module DIGITAL_CLOCK(
	RESETN, CLK,
	KEY,
   LCD_E, LCD_RS, LCD_RW,
	LCD_DATA, PIEZO
);

input RESETN, CLK;
input [4:0] KEY;
output wire LCD_E, LCD_RS, LCD_RW, PIEZO;
output wire [7:0] LCD_DATA;

wire [16:0] ALARM_TIME = 0;
wire [16:0] SETTING_TIME = 0;
wire [16:0] SETTING_DATE = 0;

wire [16:0] DISPLAY_TIME = 0;
wire [16:0] DISPLAY_DATE = 0;

wire [1:0] MODE;
wire [2:0] FLAG, CONT;

wire IS_SAVED_TIME;
wire ALARM_SET, ALARM_DOING;

// Key Controller
KEY_CONT(
	RESETN, CLK,
	KEY, DISPLAY_TIME,
	MODE, FLAG, CONT, UP, DOWN,
	DISPLAY_TIME, SET_ALARM
);

/// Time Controller
TIME_CONT CURRENT_TIME_CONT(
	RESETN, CLK,
	DISPLAY_TIME, DISPLAY_DATE,
	FLAG, UP, DOWN,
	SETTING_TIME, SETTING_DATE
);

/// Alarm Controller
ALARM_TIME_CONT ALARM_TIME_CONT(
	RESETN, CLK,
	DISPLAY_TIME,
	FLAG, UP, DOWN,
	ALARM_TIME
);

/// Current Time Calculator
TIME_CAL CURRENT_TIME_CAL(
	RESETN, CLK,
	SETTING_TIME, SETTING_DATE, ALARM_TIME,
	IS_SAVED_TIME, FLAG,
	DISPLAY_TIME, DISPLAY_DATE
);

/// (current time) and alarm time) compare
TIME_COMPARE(
	RESETN, CLK,
	ALARM_SET, DISPLAY_TIME, ALARM_TIME,
	ALARM_DOING
);

/// PIEZO
PIEZO_UNIT(
	RESETN, CLK,
	ALARM_DOING,
	PIEZO
);

/// LCD Controller
LCD_CONT(
    RESETN, CLK,
	 DISPLAY_TIME, DISPLAY_DATE,
	 MODE, CONT, RING_ALARM, SET_ALARM,
    LCD_E, LCD_RS, LCD_RW,
    LCD_DATA
);


endmodule
