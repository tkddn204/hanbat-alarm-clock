
/* CURRENT_TIME BIT LIST
`define   IN_MERIDIAN IN_TIME[17]
`define	 IN_HOUR     IN_TIME[16:12]
`define	 IN_MIN      IN_TIME[11:6]
`define   IN_SEC      IN_TIME[5:0]

/* CURRENT_DATE BIT LIST
`define   IN_YEAR     IN_DATE[15:9]
`define	 IN_MONTH    IN_DATE[8:5]
`define	 IN_DAY      IN_DATE[4:0]
*/

/* ALARM_TIME BIT LIST
`define	 IN_HOUR     IN_TIME[16:12]
`define	 IN_MIN      IN_TIME[11:6]
`define   IN_SEC      IN_TIME[5:0]
*/

// DISPLAY_CONT.v

module DISPLAY_CONT(
	RESETN, CLK,
	CURRENT_TIME, CURRENT_DATE, ALARM_TIME,
	MODE, ALARM_ENABLE, ALARM_DOING,
	DISPLAY_DATA
);

input RESETN, CLK;
input [4:0] KEY;
input [16:0] ALARM_TIME;
input [17:0] CURRENT_TIME;
input [15:0] CURRENT_DATE;
input [5:0] MODE;
input ALARM_ENABLE, ALARM_DOING;
// LINE 1 -> [15:0], LINE 2 -> [31:16]
input [7:0] DISPLAY_DATA [31:0];

wire [7:0] H10, H1, M10, M1, S10, S1, M;
wire [7:0] Y10, Y1, MT10, MT1, D10, D1;

wire [7:0] OUT_H10, OUT_H1, OUT_M10, OUT_M1, OUT_S10, OUT_S1;
wire [7:0] OUT_Y10, OUT_Y1, OUT_MT10, OUT_MT1, OUT_D10, OUT_D1;

/* MODE */
parameter CURRENT_TIME = 6'b000000,
			 CURRENT_CONTROL_TIME = 6'b010000,
			 CURRENT_CONTROL_HOUR = 6'b010011,
			 CURRENT_CONTROL_MIN = 6'b010101,
			 CURRENT_CONTROL_SEC = 6'b010111,
			 CURRENT_CONTROL_MERIDIAN = 6'b011001,
			 CURRENT_CONTROL_YEAR = 6'b011011,
			 CURRENT_CONTROL_MONTH = 6'b011101,
			 CURRENT_CONTROL_DAY = 6'b011111,
			 ALARM_TIME = 6'b100001,
			 ALARM_CONTROL_TIME = 6'b110001,
			 ALARM_CONTROL_HOUR = 6'b110011,
			 ALARM_CONTROL_MIN = 6'b110101,
			 ALARM_CONTROL_SEC = 6'b110111;
			 
/* MERIDIAN LIST(A, B) */
parameter AM = 8'b01000001,
			 PM = 8'b01000010;
			 
// x, y, z => input x, output y, z
WT_SEP HOUR_SEP(HOUR, H10, H1);
WT_SEP MIN_SEP(MIN, M10, M1);
WT_SEP SECOND_SEP(SEC, S10, S1);

WT_SEP YEAR_SEP(YEAR, Y10, Y1);
WT_SEP MONTH_SEP(MONTH, MT10, MT1);
WT_SEP DAY_SEP(DAY, D10, D1);

// decode x to y
WT_DECODER H10_DECODE(H10, OUT_H10);
WT_DECODER H1_DECODE(H1, OUT_H1);
WT_DECODER M10_DECODE(M10, OUT_M10);
WT_DECODER M1_DECODE(M1, OUT_M1);
WT_DECODER S10_DECODE(S10, OUT_S10);
WT_DECODER S1_DECODE(S1, OUT_S1);

WT_DECODER Y10_DECODE(Y10, OUT_Y10);
WT_DECODER Y1_DECODE(Y1, OUT_Y1);
WT_DECODER MT10_DECODE(D10, OUT_MT10);
WT_DECODER MT1_DECODE(D1, OUT_MT1);
WT_DECODER D10_DECODE(D10, OUT_D10);
WT_DECODER D1_DECODE(D1, OUT_D1);

always @(posedge CLK)
begin
	if(!RESETN)
		begin
			for(integer i = 0; i < 32; i = i++)
				begin
					DISPLAY_DATA[i] = 8'b00100000;
				end
		end
	else
		begin
			
		end
end

endmodule
