module DISPLAY_DECODER(
	RESETN, CLK,
	IN_TIME, IN_DATE, IN_ALARM_TIME,
	OUT_H10, OUT_H1, OUT_M10, OUT_M1, OUT_S10, OUT_S1, OUT_MERIDIAN,
	OUT_Y10, OUT_Y1, OUT_MT10, OUT_MT1, OUT_D10, OUT_D1,
	OUT_ALARM_H10, OUT_ALARM_H1, OUT_ALARM_M10, OUT_ALARM_M1, OUT_ALARM_S10, OUT_ALARM_S1
);

input RESETN, CLK;
input [16:0] IN_ALARM_TIME;
input [17:0] IN_TIME;
input [15:0] IN_DATE;
output wire [7:0] OUT_ALARM_H10, OUT_ALARM_H1, OUT_ALARM_M10, OUT_ALARM_M1, OUT_ALARM_S10, OUT_ALARM_S1;
output wire [7:0] OUT_H10, OUT_H1, OUT_M10, OUT_M1, OUT_S10, OUT_S1, OUT_MERIDIAN;
output wire [7:0] OUT_Y10, OUT_Y1, OUT_MT10, OUT_MT1, OUT_D10, OUT_D1;

// Current
reg MERIDIAN;
reg [4:0] HOUR;
reg [5:0] MIN, SEC;

reg [6:0] YEAR;
reg [3:0] MONTH;
reg [4:0] DAY;

wire [7:0] H10, H1, M10, M1, S10, S1;
wire [7:0] Y10, Y1, MT10, MT1, D10, D1;
wire [7:0] ALARM_H10, ALARM_H1, ALARM_M10, ALARM_M1, ALARM_S10, ALARM_S1;

// Alarm
reg [4:0] ALARM_HOUR;
reg [5:0] ALARM_MIN, ALARM_SEC;

always @(posedge CLK)
begin
	if(!RESETN)
		begin
			MERIDIAN = 0;
			HOUR = 0;
			MIN  = 0;
			SEC  = 0;
			
			YEAR  = 16;
			MONTH = 1;
			DAY   = 1;
			
			ALARM_HOUR = 0;
			ALARM_MIN  = 0;
			ALARM_SEC  = 0;
		end
	else
		begin
			MERIDIAN = IN_TIME[17];
			HOUR = IN_TIME[16:12];
			MIN  = IN_TIME[11:6];
			SEC  = IN_TIME[5:0];
			
			YEAR  = IN_DATE[15:9];
			MONTH = IN_DATE[8:5];
			DAY   = IN_DATE[4:0];
			
			ALARM_HOUR = IN_ALARM_TIME[16:12];
			ALARM_MIN  = IN_ALARM_TIME[11:6];
			ALARM_SEC  = IN_ALARM_TIME[5:0];
		end
end

assign OUT_MERIDIAN = MERIDIAN;

// x, y, z => input x, output y, z
WT_SEP HOUR_SEP(HOUR, H10, H1);
WT_SEP MIN_SEP(MIN, M10, M1);
WT_SEP SECOND_SEP(SEC, S10, S1);

WT_SEP YEAR_SEP(YEAR, Y10, Y1);
WT_SEP MONTH_SEP(MONTH, MT10, MT1);
WT_SEP DAY_SEP(DAY, D10, D1);

WT_SEP ALARM_HOUR_SEP(ALARM_HOUR, ALARM_H10, ALARM_H1);
WT_SEP ALARM_MIN_SEP(ALARM_MIN, ALARM_M10, ALARM_M1);
WT_SEP ALARM_SECOND_SEP(ALARM_SEC, ALARM_S10, ALARM_S1);

// decode x to y
WT_DECODER H10_DECODE(H10, OUT_H10);
WT_DECODER H1_DECODE(H1, OUT_H1);
WT_DECODER M10_DECODE(M10, OUT_M10);
WT_DECODER M1_DECODE(M1, OUT_M1);
WT_DECODER S10_DECODE(S10, OUT_S10);
WT_DECODER S1_DECODE(S1, OUT_S1);

WT_DECODER Y10_DECODE(Y10, OUT_Y10);
WT_DECODER Y1_DECODE(Y1, OUT_Y1);
WT_DECODER MT10_DECODE(D10, OUT_MT10);
WT_DECODER MT1_DECODE(D1, OUT_MT1);
WT_DECODER D10_DECODE(D10, OUT_D10);
WT_DECODER D1_DECODE(D1, OUT_D1);

WT_DECODER ALARM_H10_DECODE(ALARM_H10, OUT_ALARM_H10);
WT_DECODER ALARM_H1_DECODE(ALARM_H1, OUT_ALARM_H1);
WT_DECODER ALARM_M10_DECODE(ALARM_M10, OUT_ALARM_M10);
WT_DECODER ALARM_M1_DECODE(ALARM_M1, OUT_ALARM_M1);
WT_DECODER ALARM_S10_DECODE(ALARM_S10, OUT_ALARM_S10);
WT_DECODER ALARM_S1_DECODE(ALARM_S1, OUT_ALARM_S1);

endmodule
